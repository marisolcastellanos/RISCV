module adder(input  [31:0] a, b,
             output [31:0] y);

  //add a to b
  
endmodule
